LIBRARY IEEE;
USE IEEE.sTD_LOGIC_1164.ALL;

PACKAGE lab3_package IS
	COMPONENT fullAdd
		PORT (
			Cin, x, y : IN STD_LOGIC;
			s, Cout : OUT STD_LOGIC
		);
	END COMPONENT fullAdd;

	COMPONENT hex
		PORT (
			I : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			O : OUT STD_LOGIC_VECTOR(0 TO 6)
		);
	END COMPONENT hex;

	COMPONENT FA4
		PORT (
			Cin : IN STD_LOGIC;
			A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			Cout : OUT STD_LOGIC
		);
	END COMPONENT FA4;

	COMPONENT BCD
		PORT (
			Cin : IN STD_LOGIC;
			A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			Cout : OUT STD_LOGIC
		);
	END COMPONENT BCD;
END lab3_package;